`timescale 1ns / 1ps

module Hamming_Decoder(
    input wire [6:0] IN,
    input wire CLK, 
    input wire RESET,
    output wire [3:0] OUT
);




endmodule

